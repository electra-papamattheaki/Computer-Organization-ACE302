----------------------------------------------------------------------------------
-- Decoder 5-to-32.
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Decoder is
    Port ( decoder_in : in STD_LOGIC_VECTOR (4 downto 0);
           decoder_out : out STD_LOGIC_VECTOR (31 downto 0));
end Decoder;

architecture Behavioral_Decoder of Decoder is

begin
    
    -- Using HEX Form for the output to make it easier for the simulation
    with (decoder_in) select
        decoder_out <= X"00000001" when "00000", -- 0
                       X"00000002" when "00001", -- 1
                       X"00000004" when "00010", -- 2
                       X"00000008" when "00011", -- 3
                       X"00000010" when "00100", -- 4
                       X"00000020" when "00101", -- 5
                       X"00000040" when "00110", -- 6
                       X"00000080" when "00111", -- 7
                       X"00000100" when "01000", -- 8
                       X"00000200" when "01001", -- 9
                       X"00000400" when "01010", -- 10
                       X"00000800" when "01011", -- 11
                       X"00001000" when "01100", -- 12
                       X"00002000" when "01101", -- 13
                       X"00004000" when "01110", -- 14
                       X"00008000" when "01111", -- 15
                       X"00010000" when "10000", -- 16
                       X"00020000" when "10001", -- 17
                       X"00040000" when "10010", -- 18
                       X"00080000" when "10011", -- 19
                       X"00100000" when "10100", -- 20
                       X"00200000" when "10101", -- 21
                       X"00400000" when "10110", -- 22
                       X"00800000" when "10111", -- 23
                       X"01000000" when "11000", -- 24
                       X"02000000" when "11001", -- 25
                       X"04000000" when "11010", -- 26
                       X"08000000" when "11011", -- 27
                       X"10000000" when "11100", -- 28
                       X"20000000" when "11101", -- 29
                       X"40000000" when "11110", -- 30
                       X"80000000" when "11111", -- 31
                       X"00000000" when others;  -- all off
                       
--  Another way using 32-bit form for the output
--        with (decoder_in) select
--        decoder_out <= "00000000000000000000000000000001" when "00000", -- 0
--                       "00000000000000000000000000000010" when "00001", -- 1
--                       "00000000000000000000000000000100" when "00010", -- 2
--                       "00000000000000000000000000001000" when "00011", -- 3
--                       "00000000000000000000000000010000" when "00100", -- 4
--                       "00000000000000000000000000100000" when "00101", -- 5
--                       "00000000000000000000000001000000" when "00110", -- 6
--                       "00000000000000000000000010000000" when "00111", -- 7
--                       "00000000000000000000000100000000" when "01000", -- 8
--                       "00000000000000000000001000000000" when "01001", -- 9
--                       "00000000000000000000010000000000" when "01010", -- 10
--                       "00000000000000000000100000000000" when "01011", -- 11
--                       "00000000000000000001000000000000" when "01100", -- 12
--                       "00000000000000000010000000000000" when "01101", -- 13
--                       "00000000000000000100000000000000" when "01110", -- 14
--                       "00000000000000010000000000000000" when "01111", -- 15
--                       "00000000000000100000000000000000" when "10000", -- 16
--                       "00000000000001000000000000000000" when "10001", -- 17
--                       "00000000000010000000000000000000" when "10010", -- 18
--                       "00000000000100000000000000000000" when "10011", -- 19
--                       "00000000001000000000000000000000" when "10100", -- 20
--                       "00000000010000000000000000000000" when "10101", -- 21
--                       "00000000100000000000000000000000" when "10110", -- 22
--                       "00000001000000000000000000000000" when "10111", -- 23
--                       "00000010000000000000000000000000" when "11000", -- 24
--                       "00000100000000000000000000000000" when "11001", -- 25
--                       "00001000000000000000000000000000" when "11010", -- 26
--                       "00010000000000000000000000000000" when "11011", -- 27
--                       "00010000000000000000000000000000" when "11100", -- 28
--                       "00100000000000000000000000000000" when "11101", -- 29
--                       "01000000000000000000000000000000" when "11110", -- 30
--                       "10000000000000000000000000000000" when "11111"; -- 31
        
end Behavioral_Decoder;
